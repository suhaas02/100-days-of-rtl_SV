module clock_generator(clock); 
    input clock; 
    //initial clock = 0; 
    //always #10 clock = ~clock;
endmodule  